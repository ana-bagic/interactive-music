BZh91AY&SY��Ի �_�Px��g߰����P�Ӵ1��+N�R�Ҙ����M� �j0�f����(bm#d`�4�		i�7�6��zhF��  OQ�C�L`�a4� d�@�E4��{�S�M��h i�2����I] 4 PI��$:�i.I��M��!X0Tb�5&MX��9���ǲ�������u��㲝.V���}�e0 �̮��uQG:��sz���U�.v���´��Neq?H�h�Lf�����s��Ů[:���DDDa�Zh�cL|.�٢���Υ�T����s&#��56�(b*��2������;�'@�x�Li����x�|�2�c.SaP��yJ�S�U$�N+WB�֎3���z��TY���Z�_)��H�j��驹Ą&6�m�An��/��(���NkH�LC09lC����2��%S),YI��u�Dj�e�8F l�3t����\�����.��ベ��aK�AWK��%�E��X�(�6��H�OtS]^D�A��P~�
�h� �h��d(��B#�ˍ~�Qx�揖�A�˥�,��!\i���yqrt���"B^�c���5m�� \�62�["C�"�,��]��َ�n�4�4s�"	�®[�����|Vb
�	�DtoGd��LW�.bۦ�K<Y��k�_��F
)њ�8��Q���b�uO5ȘZd�,�S�:Ÿ��9����@���b��]9�O:�-`J�@�_d�P2�c�?l��g(�pRRj�IRA%0{z���<���@��O((?I�v�i$�,���K3Ec��������L@�H�1���@^Rd-��
�Seh��q{��c�5��U�)i�)��z��;H<d�؃!��P6�Յ[�tl�$4wBxlC��5kA��Sa��MY�%�Φ�%U}��4�0h-�����)�tn��