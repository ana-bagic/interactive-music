BZh91AY&SY�� =߀Py��g߰����P^wu�v����	$T�<Q�jz��I�6I��i���y6�B��@      �MU��1 h��  i��&�&	��0`��$H&�����3M"=5�z5SA���i1�}B���$"�������Ɂ6��2��pHX����Q�6�nKw$�I$�I$�.�:(�����BL�%0�5�����K�"I�2�_u��	��y_p��q,}�8��X�V���WA�@��\ ��#@/�`G��؝�˂I$�K0��Ƙ��g�ު�n�٭;a2�P�kt9��ozb� U��0eČ/,�U\�������T*��ՀB��qaR�b���i2-�������
a0$ ����n��Չ���%1XR�UXP�HY�#,E*�i:+������S����we��	;k�Ъ)�By.�@�� N�/}]�z��������9DRS\na8�l/�n������
1Q�L�j��>|^���O�#��֯ik�óN�#��������f<�\6W�]<%���n�Ǩ1���4���ا,�|��>��E��(J��G��6�A�8F�#��μ�Q���G�"��:`ы#��Uv��x]i���)Jخ㫑O~nP�
Ho�h>���h7�Pt�i�"���2ף���e�`�CC�ڨO���`��ma�q�4���C�c~�`d	�N[��f����S)��a�h6?^���#�H�3�GMt�؁_�c���Xt��Ʌ�h�wO��K�i�-PE�M���I#��3��,��@`�
{s 		������02VRu��5'�9̬5HNP�էlCVx�\Ź���{�� ��[ֳ�]<�yW�6�Z���j0��!<7�5��j�H��.tn��ȣd�ጷ�Yg�(�R��N��I�e����-K����h35��8{12C��Pת�7:CG�H0�$?̂�w�+ʬm�W
�˷$Y��ED�Zn�Z/����)����