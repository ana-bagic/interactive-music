BZh91AY&SY	��� �_�Px��g߰����P�wmcv���I�G�M��mS�4h=M  �A��	SM454���     �)5L��z���� yF� ��&0a0�` 2i�a"AOF�6)蘘2 4i|Ї���I%D���'��x0&�]�C]�t��i
т�3P��V�/!��m�d��IV��I�S�'�[b����:FB�D�.�+_J}���q�O!F�`�W��g����|��q���HE*c!���;�����X�I'&�A��B�.9u}[��L8�'�����61��$F��:�.�K^`����`!d4�+LJ�)aaUzM\%BH��Y�@vE!L.RTK�u�¶��Zԓ�r�ֹ�'PB�V�qr_�8d��,1�Y�W`���AIjI$�c:{��a��:��%�>�l$V�� ���[�)�:�L�JCZ���^��R�"�*�t��}/���F.�a����w����9l�OJ�l�cV�z3���Xcz%T�(3����Yz�\��L�Р��&7Z�R����:��%�1��`��[Af(��2b���ނ��]6����ͤDJV��7rU�f�C�����ܪ�m)ڝitd?�-�����9 i�q���O���B�~܃�A5B\�����."I�ݶ���&HݕA�A���Qy�H�$k�Aoy��^i@]���xb�'�lL.4�KJ�|g(���;�g���qSQ&,䑚s�Oo�%s )㜀$�u��yZ�Vp�Y"�T�(�B�=}��� 8��q�?L�����^��VLW�#d
y ��	3{X[1�#rc^UѾ��+2KZ6�Y�$aC6d@�R���Ǟ����^U���kL��J�( �h�D���!�0bzP)�y��HCG��a�?a� ��WB��������F�y�Rϕ���٬���"�(H��S 