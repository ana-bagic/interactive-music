BZh91AY&SY�<� #�_�Ry����߰����`�|�,�� ��z*�� � H  	  	  x���٪������Bx�d��  �~%IE�24  ���8ɓM0�14`� Ѧ z4���@      I���A����=OH4��4�# *)� &�S��G���L�h4M:��}{D�)�BO�SL�h��	�˹�T@0����_���v���Pj"$��qO���� e&�42�	.-��fI*I�(9��,��������h�^��g�������p�9ÂtzgF[��~(K%�j-�l-�d�B�[��-al-B�-E��-��Z�j�E��E��Z�աlKB@$Y$X̺}8	��3V�
��7�(��
!l+��o�3s=����;vnk]�P��RP�D�����<Q���½Y����2`�[�� ��-i*�V[nɵ[1��P@���t���9X�����b��`���i�Q�VV\�EN�mY�(���#�̏�w�AWg,�����,<cFj��[g�-�ʫ�t�#7m��N�q\�o���+>�],	Ti7Nl��A�6�(��d췒G.����� �B��yK+&�T�˕X68^�ͦ�@S��k�l�jn�Q�ȑ�:�iב���]�Hg��Ҧ������Y;AB�L]��u҆�\�(2�A�ڳ�c��2�	�@�ӦJ5č�:�T1P�� duU`�E�vH6'rB�T[pN"��BY+��&�V�j$��HƪR�A���U��T!*u��Qׄ��+@ԍ�buDd2�����M��SPn9E](���X�pr� rX2IF��&D+rU$vKF��-uR�\���H\jY��FT�VT�%L�Ue���9d��S�E��k���	$�\��� �ߏ>\������2j���C�C����-�Q_�S��@"Da;�����liq<��|όļ5�H����O��J��ѱ�rX�S�*:� �uڝn�b���؊LY�3]�|[����E$j9����w��"ĸ1$�lڲ���k,FT�W&�k�}�eL�5��&�q���(֡£joM� �gdbC��u�*�L6����d3�C�`�O�~���vn��X�yȲ���Js��ts�TTçЩ���΅ƚb͐.Zf&�W� �,�ܚ�Ng"�2��s�7.�mjѼw/�! ��{�t�!��4�P@M��x�� b�iM�y�P�O������.��B�S�d/D5�S)��pO0�'S,���}v��u¬�<�c�6��]�~�W��BBʹuBƼ���j�k��o�J��)H�G���>j�R�L/���"6�ךsg
-�v�u�=���:߱����٥?iDB� -.*q�;�[0��2t|5bU�3���4�Y��m<g��k��}�tĜ���2�����~̂~�o�5��y��o��H�֝����W�x�S��]b��Å�ڡ��ƾ/�ݩ$�4�9�BG�t�%^��we����5ޱy˘�'���>������~nb�_�{�ݎ��ʲ2��xf�© ��]�[@���޲_	������.�*������g"����Ĝ��:��(�Te��l���CG?a�{4��aE���WsE��k{��[��,���;��
�$�O~ά�`�=��A�%\��Ƽn���m�r�Ϸ���iY\F���'��l
�)y�
H��W�<��c�?�E�O�����
$��W�g9��YѲ~P��!v#��+�̵�Ŗ�n~%3vlW���A��׵���>�b�)Tf6�i��+�m�%�!TqQ�F��KN&
B�2��)X1�����܏�U Y��x~y��Zo��y�B�M��U�.��M��/�z����՚�/0�p.����X$AO�-���j������0�wX���#�ckDKQ�1����&����j����O�#dt2D�GΠ���y�R��
|����ϱ3���sKq�*>��x��c�����F}ળh�*v�|sm���5��ޕP�n�
D?&����]�wW�F�j��#
�x/9jsg�dL묠Sʻ��ѨoN�v�m8��*e\��c��6µ������&*��[�0x�%�0�3T2�7������S:�NvEc3��v.���l�}{[�x�/�[���v����D̶�*$��B�Br�r˼����M��߹a{~:��	Y�rJ�\]���Q�� l7+K���Mo�:m�w-I^��!���{��Iy�s�%Zo�+�4=��NM��^QI�L)�
��k�h{�_5b]͋J��W� ���UCT��Tŕ����u}��R6�_>y�E�M�Ī��׻�-{�0鷘�g+!%C+w��o�`�P�|%��5��>o���W���ug'oQ�y��RD�nO]�t�#pR���qQT�]��T9$dhp�8Q���(���m�։*7LQ����jʅ�Nb���ig�W[�t7_�Ei�`�Fj�4b�?:��ޛ��W��7+o��k}�M�Xr�R��>���y���ۻ�x��-^����YR�C ���'��g-�'!V���fw��]B�إ�	����x�Υ��'�G�~�3k0�������ƭ�,�n*该�5Xs�pF�#VꇏaU��q����$�Q��z�Q`��rm�D�v���,Y�Խ�oA����)��ܱE�M�&43��3߷�����;�B���n᫆���wq�y)<?F����g����n���Z�ƗX��"�<0vmZ�4��4�3������(��1v��V��	�LFik�ۋ��޿Qг/��$-ȖP��ׁ��w��K�l��ii�ؼoÎ���瓫O ��I#i��7k'U�喍jU�mcU�����Un��y��&\��B�?vF`��(��\k؄~����J��ƍ���aE��5?�Ŷw�j�_h�ݹ��Ԇ1Q_:�F c�4��[YR�VJ�j
Yk��$d�;j���Ԓ����5���`���C���r����+�o���%���i�[ʏ����yU��=���vn��S�G�Z=WjB|5$s�ڣR�]��7>��m�J\�˿rR�o�LK[罴����񺺩Bs<5h�1z�b�S��U�M�/vU/|��h��Ij4JE��L<������Ӓ�}���M�Vfp�\�=����S�.��={���]�v�(�S�f{�}{ޢI��v#���O�z�%��"W���G��τ����Hm��o�Tݮ������Q�jm��Gh����w��O��֔�%��e�S||�=J��߳��"x��ǔ�h�uoɣ�H6�*����ƞ��(���t=�z+�3�uo��з�8I ��d�{Լ�^ط:��Q�� W�U�]ߠل�-4�^U�8����G��/UU��˧N�T�X˝�	������c3m�Ddm�#uWe �jI-hj��ZSCg��nj�*����n{�F����������u��٫	�tܠl���|}�z]
��W���_�.�'��o{��Ү��/��¿71V��ׅ#~�"�b5m�az��^Ml��sW��������4����T$��3�[��)�`�C�0��=�	�\�3�7�����yxF/��"l��{4�4.WJ�2]8�����o���e����V�����xT���-���9�{�aλ�iΜ���˭�qz��U����>�l���v��>K~�����@Tm�|+���	U�ܮH�tZk���w=*Ա����9U����%ˆ�aL3ׇ8��a���v�d�3r�%ŲF#a��r����~<�תo�r�*��K���)����g��G�fj³�$��[z�������4#��˶��%�"�e0�G?�<F��9�;N4�!D��$���FA"�D���T��o8
�>�$�3=+bҴ�Դ�����u
.���ʴ�G��@��V�kt,Vb��H�1��b)�R����-��aE�BФ�DA��7T.D�Q$�ay
�%�T)Z��B�4޲3� !h����
ʦ9��Vlni�qMf�g��]K���I$Z	-��Ŷ�����X�|��Y�N��7c� l�#磆��A�{��G��kn�erݿ�{cQ�g����=��oo<� �}������|\�gzE9�&ga����&:��*�^D�?[\ؖ��x�1.���5Mj���a����t�������v]}�� ��)���x�!Bl��{i�!�`����h��O�24C���~飏����?��:�9��8>�|�c꾏*���p����|4�I���4����Qb�R�L�?`�����RLi�f��(�a������!�<(�p��RE��my%��0��G݉i�+�4�
بF����d1H�� ����Q1�1+GLpQ�LL�m�ђ}MN�i���r\�PWXRh�H��m���ޖ7������B�g��ӌ؛�9���B7�z��n��W�����<<�V
�$��L\����\��p���v;6d�f���7'V\[H�,���8'qy{ڞ�Y=§�ָ�<�s
���:y��Ν[�¨m�!6��X�^��sc�	���>)Ot�b�"��ࢁ��yU�����B#���O�X��0��C��N1�ٹ���,#�1WΆ�A�0r�#�Xi�l)c���ږ�PP/eq㠸��|�6+���]Y&��D���Z��bT�#�y��lNCI.��d�,2�4��k�m�e6�n���%{|�������$@��|_X}
�;�߮}�*O����:�OWN��9p�����%�6
�v<����{[�=f�/��N��m�.�Qq:g�~�b�f�F��|��r{�xe��{��4����896� ��p�l~'.C��M�*]P�t�{�#�%щ10�X�"Hb��4�ݭ�e��/�g !���R���@�b`�P�l	��/7	"ǎc���v8ip���j�"�'<%��#��p�lvDṹ��n���S$1$����������1yB��
n�jʄr�'�����:�d����wF����w����P��E)�u:5D���m �8QH����#��b9����)�t��